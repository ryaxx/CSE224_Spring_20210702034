VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO my_first_design
  CLASS BLOCK ;
  FOREIGN my_first_design ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 50.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.020 10.640 39.620 38.320 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.380 44.400 19.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 10.640 36.320 38.320 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.080 44.400 16.680 ;
    END
  END VPWR
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END in[0]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END in[7]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 43.560 50.000 44.160 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 38.120 50.000 38.720 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 32.680 50.000 33.280 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 27.240 50.000 27.840 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 21.800 50.000 22.400 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 16.360 50.000 16.960 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 10.920 50.000 11.520 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 5.480 50.000 6.080 ;
    END
  END out[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 44.350 38.165 ;
      LAYER li1 ;
        RECT 5.520 10.795 44.160 38.165 ;
      LAYER met1 ;
        RECT 4.210 10.640 44.160 38.320 ;
      LAYER met2 ;
        RECT 4.230 5.595 42.230 44.045 ;
      LAYER met3 ;
        RECT 4.400 43.160 45.600 44.025 ;
        RECT 3.990 39.120 46.000 43.160 ;
        RECT 4.400 37.720 45.600 39.120 ;
        RECT 3.990 33.680 46.000 37.720 ;
        RECT 4.400 32.280 45.600 33.680 ;
        RECT 3.990 28.240 46.000 32.280 ;
        RECT 4.400 26.840 45.600 28.240 ;
        RECT 3.990 22.800 46.000 26.840 ;
        RECT 4.400 21.400 45.600 22.800 ;
        RECT 3.990 17.360 46.000 21.400 ;
        RECT 4.400 15.960 45.600 17.360 ;
        RECT 3.990 11.920 46.000 15.960 ;
        RECT 4.400 10.520 45.600 11.920 ;
        RECT 3.990 6.480 46.000 10.520 ;
        RECT 4.400 5.615 45.600 6.480 ;
  END
END my_first_design
END LIBRARY

