magic
tech sky130A
magscale 1 2
timestamp 1745779526
<< nwell >>
rect 1066 2159 8870 7633
<< obsli1 >>
rect 1104 2159 8832 7633
<< obsm1 >>
rect 842 2128 8832 7664
<< obsm2 >>
rect 846 1119 8446 8809
<< metal3 >>
rect 0 8712 800 8832
rect 9200 8712 10000 8832
rect 0 7624 800 7744
rect 9200 7624 10000 7744
rect 0 6536 800 6656
rect 9200 6536 10000 6656
rect 0 5448 800 5568
rect 9200 5448 10000 5568
rect 0 4360 800 4480
rect 9200 4360 10000 4480
rect 0 3272 800 3392
rect 9200 3272 10000 3392
rect 0 2184 800 2304
rect 9200 2184 10000 2304
rect 0 1096 800 1216
rect 9200 1096 10000 1216
<< obsm3 >>
rect 880 8632 9120 8805
rect 798 7824 9200 8632
rect 880 7544 9120 7824
rect 798 6736 9200 7544
rect 880 6456 9120 6736
rect 798 5648 9200 6456
rect 880 5368 9120 5648
rect 798 4560 9200 5368
rect 880 4280 9120 4560
rect 798 3472 9200 4280
rect 880 3192 9120 3472
rect 798 2384 9200 3192
rect 880 2104 9120 2384
rect 798 1296 9200 2104
rect 880 1123 9120 1296
<< metal4 >>
rect 1944 2128 2264 7664
rect 2604 2128 2924 7664
rect 6944 2128 7264 7664
rect 7604 2128 7924 7664
<< metal5 >>
rect 1056 3676 8880 3996
rect 1056 3016 8880 3336
<< labels >>
rlabel metal4 s 2604 2128 2924 7664 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 7664 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3676 8880 3996 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3016 8880 3336 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 8712 800 8832 6 in[0]
port 3 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 in[1]
port 4 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 in[2]
port 5 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 in[3]
port 6 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 in[4]
port 7 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 in[5]
port 8 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 in[6]
port 9 nsew signal input
rlabel metal3 s 0 1096 800 1216 6 in[7]
port 10 nsew signal input
rlabel metal3 s 9200 8712 10000 8832 6 out[0]
port 11 nsew signal output
rlabel metal3 s 9200 7624 10000 7744 6 out[1]
port 12 nsew signal output
rlabel metal3 s 9200 6536 10000 6656 6 out[2]
port 13 nsew signal output
rlabel metal3 s 9200 5448 10000 5568 6 out[3]
port 14 nsew signal output
rlabel metal3 s 9200 4360 10000 4480 6 out[4]
port 15 nsew signal output
rlabel metal3 s 9200 3272 10000 3392 6 out[5]
port 16 nsew signal output
rlabel metal3 s 9200 2184 10000 2304 6 out[6]
port 17 nsew signal output
rlabel metal3 s 9200 1096 10000 1216 6 out[7]
port 18 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 200484
string GDS_FILE /openlane/designs/my_first_design/runs/RUN_2025.04.27_18.41.48/results/signoff/my_first_design.magic.gds
string GDS_START 105490
<< end >>

