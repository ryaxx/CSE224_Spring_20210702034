module InstructionMemory(input [4:0] addr, output reg [31:0] instr);
    always @(*) begin
        case(addr)
            0: instr = 32'b110_00000_01010_0000000000001010;  // ADDI r10, r0, 10
            1: instr = 32'b110_00000_01111_0000000000001111;  // ADDI r15, r0, 15
            2: instr = 32'b010_01010_01111_11001_00000000000; // ADD r25, r10, r15
            3: instr = 32'b111_11001_10100_0000000000000101;  // SUBI r20, r25, 5
            4: instr = 32'b110_00000_10101_0000000000000010;  // ADDI r21, r0, 2
            5: instr = 32'b000_00000_00000_00000_00000001100; // J 12
            12: instr = 32'b110_00000_00100_0000000000000100; // ADDI r4, r0, 4
            13: instr = 32'b010_00000_00000_00101_00000000000; // ADD r5, r0, r0
            14: instr = 32'b001_00100_00101_00000_00000000111; // BEQ r4, r5, 7
            15: instr = 32'b110_00000_00110_0000000000000001; // ADDI r6, r0, 1
            16: instr = 32'b110_00000_00111_0000000000000001; // ADDI r7, r0, 1
            17: instr = 32'b010_00110_00111_01000_00000000000; // ADD r8, r6, r7
            18: instr = 32'b010_00111_00000_00110_00000000000; // ADD r6, r7, r0
            19: instr = 32'b010_01000_00000_00111_00000000000; // ADD r7, r8, r0
            20: instr = 32'b110_00101_00101_0000000000000001; // ADDI r5, r5, 1
            21: instr = 32'b000_00000_00000_00000_00000001110; // J 14
            default: instr = 32'b0;
        endcase
    end
endmodule

