magic
tech sky130A
magscale 1 2
timestamp 1745779542
<< checkpaint >>
rect -3932 -2836 13932 12764
<< viali >>
rect 8033 7497 8067 7531
rect 8401 7497 8435 7531
rect 1409 7361 1443 7395
rect 3985 7361 4019 7395
rect 7849 7361 7883 7395
rect 8217 7361 8251 7395
rect 1685 7293 1719 7327
rect 3893 7293 3927 7327
rect 4353 7157 4387 7191
rect 1501 6749 1535 6783
rect 1777 6749 1811 6783
rect 2053 6749 2087 6783
rect 6101 6749 6135 6783
rect 6285 6749 6319 6783
rect 7205 6749 7239 6783
rect 7389 6749 7423 6783
rect 8217 6749 8251 6783
rect 1593 6613 1627 6647
rect 1961 6613 1995 6647
rect 2237 6613 2271 6647
rect 6469 6613 6503 6647
rect 7297 6613 7331 6647
rect 8401 6613 8435 6647
rect 2329 6409 2363 6443
rect 6561 6341 6595 6375
rect 2145 6273 2179 6307
rect 6469 6273 6503 6307
rect 1961 6205 1995 6239
rect 6929 6205 6963 6239
rect 6745 6069 6779 6103
rect 7849 5865 7883 5899
rect 2421 5797 2455 5831
rect 5365 5729 5399 5763
rect 7389 5729 7423 5763
rect 1409 5661 1443 5695
rect 2237 5661 2271 5695
rect 2421 5661 2455 5695
rect 5457 5661 5491 5695
rect 7481 5661 7515 5695
rect 8217 5661 8251 5695
rect 1593 5525 1627 5559
rect 5825 5525 5859 5559
rect 8401 5525 8435 5559
rect 6653 5321 6687 5355
rect 2421 5185 2455 5219
rect 2697 5185 2731 5219
rect 6469 5185 6503 5219
rect 2513 5117 2547 5151
rect 2513 4981 2547 5015
rect 2881 4981 2915 5015
rect 1593 4777 1627 4811
rect 3893 4777 3927 4811
rect 4169 4777 4203 4811
rect 4169 4641 4203 4675
rect 1409 4573 1443 4607
rect 4077 4573 4111 4607
rect 8217 4573 8251 4607
rect 4353 4505 4387 4539
rect 8401 4437 8435 4471
rect 1961 4097 1995 4131
rect 2053 4097 2087 4131
rect 2237 4097 2271 4131
rect 2145 4029 2179 4063
rect 2421 3893 2455 3927
rect 1593 3689 1627 3723
rect 5733 3689 5767 3723
rect 6377 3689 6411 3723
rect 5825 3621 5859 3655
rect 6193 3553 6227 3587
rect 6285 3553 6319 3587
rect 1409 3485 1443 3519
rect 6469 3485 6503 3519
rect 6561 3485 6595 3519
rect 8217 3485 8251 3519
rect 8401 3349 8435 3383
rect 2605 3145 2639 3179
rect 2237 3009 2271 3043
rect 2329 3009 2363 3043
rect 4813 3009 4847 3043
rect 4997 2873 5031 2907
rect 2237 2805 2271 2839
rect 1593 2601 1627 2635
rect 1869 2601 1903 2635
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 7849 2397 7883 2431
rect 8217 2397 8251 2431
rect 8033 2261 8067 2295
rect 8401 2261 8435 2295
<< metal1 >>
rect 1104 7642 8832 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 8832 7642
rect 1104 7568 8832 7590
rect 8018 7488 8024 7540
rect 8076 7488 8082 7540
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 842 7352 848 7404
rect 900 7392 906 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 900 7364 1409 7392
rect 900 7352 906 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8018 7392 8024 7404
rect 7883 7364 8024 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1636 7296 1685 7324
rect 1636 7284 1642 7296
rect 1673 7293 1685 7296
rect 1719 7293 1731 7327
rect 1673 7287 1731 7293
rect 3602 7284 3608 7336
rect 3660 7324 3666 7336
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 3660 7296 3893 7324
rect 3660 7284 3666 7296
rect 3881 7293 3893 7296
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 4338 7148 4344 7200
rect 4396 7148 4402 7200
rect 1104 7098 8832 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 8832 7098
rect 1104 7024 8832 7046
rect 1486 6740 1492 6792
rect 1544 6740 1550 6792
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 934 6672 940 6724
rect 992 6712 998 6724
rect 1780 6712 1808 6743
rect 1854 6740 1860 6792
rect 1912 6740 1918 6792
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 5718 6780 5724 6792
rect 2087 6752 5724 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 6086 6740 6092 6792
rect 6144 6740 6150 6792
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 6362 6740 6368 6792
rect 6420 6780 6426 6792
rect 7193 6783 7251 6789
rect 7193 6780 7205 6783
rect 6420 6752 7205 6780
rect 6420 6740 6426 6752
rect 7193 6749 7205 6752
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 7524 6752 8217 6780
rect 7524 6740 7530 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 992 6684 1808 6712
rect 1872 6712 1900 6740
rect 1872 6684 2268 6712
rect 992 6672 998 6684
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1670 6644 1676 6656
rect 1627 6616 1676 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2240 6653 2268 6684
rect 1949 6647 2007 6653
rect 1949 6644 1961 6647
rect 1912 6616 1961 6644
rect 1912 6604 1918 6616
rect 1949 6613 1961 6616
rect 1995 6613 2007 6647
rect 1949 6607 2007 6613
rect 2225 6647 2283 6653
rect 2225 6613 2237 6647
rect 2271 6613 2283 6647
rect 2225 6607 2283 6613
rect 6454 6604 6460 6656
rect 6512 6604 6518 6656
rect 7282 6604 7288 6656
rect 7340 6604 7346 6656
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 1104 6554 8832 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 8832 6554
rect 1104 6480 8832 6502
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 7374 6440 7380 6452
rect 2363 6412 7380 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 6549 6375 6607 6381
rect 6549 6372 6561 6375
rect 4120 6344 6561 6372
rect 4120 6332 4126 6344
rect 6549 6341 6561 6344
rect 6595 6341 6607 6375
rect 6549 6335 6607 6341
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6304 2191 6307
rect 2406 6304 2412 6316
rect 2179 6276 2412 6304
rect 2179 6273 2191 6276
rect 2133 6267 2191 6273
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 6086 6264 6092 6316
rect 6144 6304 6150 6316
rect 6457 6307 6515 6313
rect 6457 6304 6469 6307
rect 6144 6276 6469 6304
rect 6144 6264 6150 6276
rect 6457 6273 6469 6276
rect 6503 6273 6515 6307
rect 6457 6267 6515 6273
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6236 2007 6239
rect 2314 6236 2320 6248
rect 1995 6208 2320 6236
rect 1995 6205 2007 6208
rect 1949 6199 2007 6205
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 3936 6208 6929 6236
rect 3936 6196 3942 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 6733 6103 6791 6109
rect 6733 6069 6745 6103
rect 6779 6100 6791 6103
rect 7558 6100 7564 6112
rect 6779 6072 7564 6100
rect 6779 6069 6791 6072
rect 6733 6063 6791 6069
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 1104 6010 8832 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 8832 6010
rect 1104 5936 8832 5958
rect 7837 5899 7895 5905
rect 7837 5865 7849 5899
rect 7883 5896 7895 5899
rect 8202 5896 8208 5908
rect 7883 5868 8208 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 2409 5831 2467 5837
rect 2409 5797 2421 5831
rect 2455 5828 2467 5831
rect 6362 5828 6368 5840
rect 2455 5800 6368 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 5368 5769 5396 5800
rect 6362 5788 6368 5800
rect 6420 5788 6426 5840
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5729 5411 5763
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 5353 5723 5411 5729
rect 5552 5732 7389 5760
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2314 5692 2320 5704
rect 2271 5664 2320 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 2406 5652 2412 5704
rect 2464 5652 2470 5704
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 2556 5664 5457 5692
rect 2556 5652 2562 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 4246 5584 4252 5636
rect 4304 5624 4310 5636
rect 5552 5624 5580 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 6546 5652 6552 5704
rect 6604 5692 6610 5704
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 6604 5664 7481 5692
rect 6604 5652 6610 5664
rect 7469 5661 7481 5664
rect 7515 5661 7527 5695
rect 7469 5655 7527 5661
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 7616 5664 8217 5692
rect 7616 5652 7622 5664
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 4304 5596 5580 5624
rect 4304 5584 4310 5596
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 4062 5556 4068 5568
rect 1627 5528 4068 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 6638 5556 6644 5568
rect 5859 5528 6644 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8389 5559 8447 5565
rect 8389 5556 8401 5559
rect 8260 5528 8401 5556
rect 8260 5516 8266 5528
rect 8389 5525 8401 5528
rect 8435 5525 8447 5559
rect 8389 5519 8447 5525
rect 1104 5466 8832 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 8832 5466
rect 1104 5392 8832 5414
rect 6641 5355 6699 5361
rect 6641 5321 6653 5355
rect 6687 5352 6699 5355
rect 7466 5352 7472 5364
rect 6687 5324 7472 5352
rect 6687 5321 6699 5324
rect 6641 5315 6699 5321
rect 7466 5312 7472 5324
rect 7524 5312 7530 5364
rect 2314 5244 2320 5296
rect 2372 5284 2378 5296
rect 2372 5256 2728 5284
rect 2372 5244 2378 5256
rect 2406 5176 2412 5228
rect 2464 5216 2470 5228
rect 2700 5225 2728 5256
rect 2685 5219 2743 5225
rect 2464 5188 2636 5216
rect 2464 5176 2470 5188
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 1636 5120 2513 5148
rect 1636 5108 1642 5120
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 2608 5148 2636 5188
rect 2685 5185 2697 5219
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 6454 5176 6460 5228
rect 6512 5176 6518 5228
rect 3878 5148 3884 5160
rect 2608 5120 3884 5148
rect 2501 5111 2559 5117
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 2498 4972 2504 5024
rect 2556 4972 2562 5024
rect 2869 5015 2927 5021
rect 2869 4981 2881 5015
rect 2915 5012 2927 5015
rect 3602 5012 3608 5024
rect 2915 4984 3608 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 1104 4922 8832 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 8832 4922
rect 1104 4848 8832 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 2314 4808 2320 4820
rect 1627 4780 2320 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 3878 4768 3884 4820
rect 3936 4768 3942 4820
rect 4154 4768 4160 4820
rect 4212 4768 4218 4820
rect 1486 4632 1492 4684
rect 1544 4672 1550 4684
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 1544 4644 4169 4672
rect 1544 4632 1550 4644
rect 4157 4641 4169 4644
rect 4203 4672 4215 4675
rect 6546 4672 6552 4684
rect 4203 4644 6552 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 7282 4564 7288 4616
rect 7340 4604 7346 4616
rect 8205 4607 8263 4613
rect 8205 4604 8217 4607
rect 7340 4576 8217 4604
rect 7340 4564 7346 4576
rect 8205 4573 8217 4576
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 4246 4496 4252 4548
rect 4304 4536 4310 4548
rect 4341 4539 4399 4545
rect 4341 4536 4353 4539
rect 4304 4508 4353 4536
rect 4304 4496 4310 4508
rect 4341 4505 4353 4508
rect 4387 4505 4399 4539
rect 4341 4499 4399 4505
rect 8386 4428 8392 4480
rect 8444 4428 8450 4480
rect 1104 4378 8832 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 8832 4378
rect 1104 4304 8832 4326
rect 2406 4196 2412 4208
rect 2056 4168 2412 4196
rect 1578 4088 1584 4140
rect 1636 4128 1642 4140
rect 2056 4137 2084 4168
rect 2406 4156 2412 4168
rect 2464 4156 2470 4208
rect 1949 4131 2007 4137
rect 1949 4128 1961 4131
rect 1636 4100 1961 4128
rect 1636 4088 1642 4100
rect 1949 4097 1961 4100
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2314 4128 2320 4140
rect 2271 4100 2320 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 2498 4060 2504 4072
rect 2179 4032 2504 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 1854 3952 1860 4004
rect 1912 3992 1918 4004
rect 2314 3992 2320 4004
rect 1912 3964 2320 3992
rect 1912 3952 1918 3964
rect 2314 3952 2320 3964
rect 2372 3992 2378 4004
rect 4154 3992 4160 4004
rect 2372 3964 4160 3992
rect 2372 3952 2378 3964
rect 4154 3952 4160 3964
rect 4212 3952 4218 4004
rect 2409 3927 2467 3933
rect 2409 3893 2421 3927
rect 2455 3924 2467 3927
rect 6178 3924 6184 3936
rect 2455 3896 6184 3924
rect 2455 3893 2467 3896
rect 2409 3887 2467 3893
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 1104 3834 8832 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 8832 3834
rect 1104 3760 8832 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 2498 3720 2504 3732
rect 1627 3692 2504 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 5718 3680 5724 3732
rect 5776 3680 5782 3732
rect 6270 3680 6276 3732
rect 6328 3720 6334 3732
rect 6365 3723 6423 3729
rect 6365 3720 6377 3723
rect 6328 3692 6377 3720
rect 6328 3680 6334 3692
rect 6365 3689 6377 3692
rect 6411 3689 6423 3723
rect 6365 3683 6423 3689
rect 3602 3612 3608 3664
rect 3660 3652 3666 3664
rect 5813 3655 5871 3661
rect 5813 3652 5825 3655
rect 3660 3624 5825 3652
rect 3660 3612 3666 3624
rect 5813 3621 5825 3624
rect 5859 3621 5871 3655
rect 5813 3615 5871 3621
rect 6178 3544 6184 3596
rect 6236 3544 6242 3596
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 842 3476 848 3528
rect 900 3516 906 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 900 3488 1409 3516
rect 900 3476 906 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 6288 3516 6316 3547
rect 4212 3488 6316 3516
rect 6457 3519 6515 3525
rect 4212 3476 4218 3488
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 4246 3408 4252 3460
rect 4304 3448 4310 3460
rect 6472 3448 6500 3479
rect 6546 3476 6552 3528
rect 6604 3476 6610 3528
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 6696 3488 8217 3516
rect 6696 3476 6702 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 4304 3420 6500 3448
rect 4304 3408 4310 3420
rect 8386 3340 8392 3392
rect 8444 3340 8450 3392
rect 1104 3290 8832 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 8832 3290
rect 1104 3216 8832 3238
rect 2593 3179 2651 3185
rect 2593 3145 2605 3179
rect 2639 3176 2651 3179
rect 6086 3176 6092 3188
rect 2639 3148 6092 3176
rect 2639 3145 2651 3148
rect 2593 3139 2651 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 4246 3108 4252 3120
rect 2240 3080 4252 3108
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 2240 3049 2268 3080
rect 4246 3068 4252 3080
rect 4304 3108 4310 3120
rect 4304 3080 4844 3108
rect 4304 3068 4310 3080
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 1728 3012 2237 3040
rect 1728 3000 1734 3012
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2314 3000 2320 3052
rect 2372 3000 2378 3052
rect 4816 3049 4844 3080
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 4985 2907 5043 2913
rect 4985 2873 4997 2907
rect 5031 2904 5043 2907
rect 8018 2904 8024 2916
rect 5031 2876 8024 2904
rect 5031 2873 5043 2876
rect 4985 2867 5043 2873
rect 8018 2864 8024 2876
rect 8076 2864 8082 2916
rect 1486 2796 1492 2848
rect 1544 2836 1550 2848
rect 2225 2839 2283 2845
rect 2225 2836 2237 2839
rect 1544 2808 2237 2836
rect 1544 2796 1550 2808
rect 2225 2805 2237 2808
rect 2271 2805 2283 2839
rect 2225 2799 2283 2805
rect 1104 2746 8832 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 8832 2746
rect 1104 2672 8832 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 3970 2632 3976 2644
rect 1903 2604 3976 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 1762 2456 1768 2508
rect 1820 2496 1826 2508
rect 1820 2468 8248 2496
rect 1820 2456 1826 2468
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 8220 2437 8248 2468
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 4396 2400 7849 2428
rect 4396 2388 4402 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8018 2252 8024 2304
rect 8076 2252 8082 2304
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 1104 2202 8832 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 8832 2202
rect 1104 2128 8832 2150
<< via1 >>
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 8024 7531 8076 7540
rect 8024 7497 8033 7531
rect 8033 7497 8067 7531
rect 8067 7497 8076 7531
rect 8024 7488 8076 7497
rect 8392 7531 8444 7540
rect 8392 7497 8401 7531
rect 8401 7497 8435 7531
rect 8435 7497 8444 7531
rect 8392 7488 8444 7497
rect 848 7352 900 7404
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 8024 7352 8076 7404
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 1584 7284 1636 7336
rect 3608 7284 3660 7336
rect 4344 7191 4396 7200
rect 4344 7157 4353 7191
rect 4353 7157 4387 7191
rect 4387 7157 4396 7191
rect 4344 7148 4396 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 1492 6783 1544 6792
rect 1492 6749 1501 6783
rect 1501 6749 1535 6783
rect 1535 6749 1544 6783
rect 1492 6740 1544 6749
rect 940 6672 992 6724
rect 1860 6740 1912 6792
rect 5724 6740 5776 6792
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6368 6740 6420 6792
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 7472 6740 7524 6792
rect 1676 6604 1728 6656
rect 1860 6604 1912 6656
rect 6460 6647 6512 6656
rect 6460 6613 6469 6647
rect 6469 6613 6503 6647
rect 6503 6613 6512 6647
rect 6460 6604 6512 6613
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 7380 6400 7432 6452
rect 4068 6332 4120 6384
rect 2412 6264 2464 6316
rect 6092 6264 6144 6316
rect 2320 6196 2372 6248
rect 3884 6196 3936 6248
rect 7564 6060 7616 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 8208 5856 8260 5908
rect 6368 5788 6420 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2320 5652 2372 5704
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 2504 5652 2556 5704
rect 4252 5584 4304 5636
rect 6552 5652 6604 5704
rect 7564 5652 7616 5704
rect 4068 5516 4120 5568
rect 6644 5516 6696 5568
rect 8208 5516 8260 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 7472 5312 7524 5364
rect 2320 5244 2372 5296
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 1584 5108 1636 5160
rect 6460 5219 6512 5228
rect 6460 5185 6469 5219
rect 6469 5185 6503 5219
rect 6503 5185 6512 5219
rect 6460 5176 6512 5185
rect 3884 5108 3936 5160
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 3608 4972 3660 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 2320 4768 2372 4820
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 4160 4811 4212 4820
rect 4160 4777 4169 4811
rect 4169 4777 4203 4811
rect 4203 4777 4212 4811
rect 4160 4768 4212 4777
rect 1492 4632 1544 4684
rect 6552 4632 6604 4684
rect 848 4564 900 4616
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 7288 4564 7340 4616
rect 4252 4496 4304 4548
rect 8392 4471 8444 4480
rect 8392 4437 8401 4471
rect 8401 4437 8435 4471
rect 8435 4437 8444 4471
rect 8392 4428 8444 4437
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 1584 4088 1636 4140
rect 2412 4156 2464 4208
rect 2320 4088 2372 4140
rect 2504 4020 2556 4072
rect 1860 3952 1912 4004
rect 2320 3952 2372 4004
rect 4160 3952 4212 4004
rect 6184 3884 6236 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 2504 3680 2556 3732
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 6276 3680 6328 3732
rect 3608 3612 3660 3664
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 848 3476 900 3528
rect 4160 3476 4212 3528
rect 4252 3408 4304 3460
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 6644 3476 6696 3528
rect 8392 3383 8444 3392
rect 8392 3349 8401 3383
rect 8401 3349 8435 3383
rect 8435 3349 8444 3383
rect 8392 3340 8444 3349
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 6092 3136 6144 3188
rect 1676 3000 1728 3052
rect 4252 3068 4304 3120
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 8024 2864 8076 2916
rect 1492 2796 1544 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 3976 2592 4028 2644
rect 1768 2456 1820 2508
rect 848 2388 900 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 4344 2388 4396 2440
rect 8024 2295 8076 2304
rect 8024 2261 8033 2295
rect 8033 2261 8067 2295
rect 8067 2261 8076 2295
rect 8024 2252 8076 2261
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
<< metal2 >>
rect 1490 8800 1546 8809
rect 1490 8735 1546 8744
rect 8022 8800 8078 8809
rect 8022 8735 8078 8744
rect 846 7576 902 7585
rect 846 7511 902 7520
rect 860 7410 888 7511
rect 848 7404 900 7410
rect 848 7346 900 7352
rect 1504 6798 1532 8735
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 8036 7546 8064 8735
rect 8390 7712 8446 7721
rect 8390 7647 8446 7656
rect 8404 7546 8432 7647
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6633 980 6666
rect 938 6624 994 6633
rect 938 6559 994 6568
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1596 5250 1624 7278
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1860 6792 1912 6798
rect 1780 6740 1860 6746
rect 1780 6734 1912 6740
rect 1780 6718 1900 6734
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1504 5222 1624 5250
rect 1504 4690 1532 5222
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 848 4616 900 4622
rect 846 4584 848 4593
rect 900 4584 902 4593
rect 846 4519 902 4528
rect 848 3528 900 3534
rect 846 3496 848 3505
rect 900 3496 902 3505
rect 846 3431 902 3440
rect 1504 2854 1532 4626
rect 1596 4146 1624 5102
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1596 2650 1624 4082
rect 1688 3058 1716 6598
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1780 2514 1808 6718
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 4010 1900 6598
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2332 5710 2360 6190
rect 2424 5710 2452 6258
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2332 5302 2360 5646
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2332 4826 2360 5238
rect 2424 5234 2452 5646
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2332 4146 2360 4762
rect 2424 4214 2452 5170
rect 2516 5030 2544 5646
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 3620 5030 3648 7278
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3896 5166 3924 6190
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2516 4078 2544 4966
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2332 3058 2360 3946
rect 2516 3738 2544 4014
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 3620 3670 3648 4966
rect 3896 4826 3924 5102
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 3988 2650 4016 7346
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4080 5574 4108 6326
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 4622 4108 5510
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4172 4010 4200 4762
rect 4264 4554 4292 5578
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4172 3534 4200 3946
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4264 3466 4292 4490
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4264 3126 4292 3402
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 1768 2508 1820 2514
rect 1768 2450 1820 2456
rect 4356 2446 4384 7142
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 5736 3738 5764 6734
rect 6104 6322 6132 6734
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 6104 3194 6132 6258
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 3602 6224 3878
rect 6288 3738 6316 6734
rect 6380 5846 6408 6734
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6472 5234 6500 6598
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6564 4690 6592 5646
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6564 3534 6592 4626
rect 6656 3534 6684 5510
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 7300 4622 7328 6598
rect 7392 6458 7420 6734
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7484 5370 7512 6734
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7576 5710 7604 6054
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 8036 2922 8064 7346
rect 8220 5914 8248 7346
rect 8392 6656 8444 6662
rect 8390 6624 8392 6633
rect 8444 6624 8446 6633
rect 8390 6559 8446 6568
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8208 5568 8260 5574
rect 8206 5536 8208 5545
rect 8260 5536 8262 5545
rect 8206 5471 8262 5480
rect 8392 4480 8444 4486
rect 8390 4448 8392 4457
rect 8444 4448 8446 4457
rect 8390 4383 8446 4392
rect 8392 3392 8444 3398
rect 8390 3360 8392 3369
rect 8444 3360 8446 3369
rect 8390 3295 8446 3304
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 1676 2440 1728 2446
rect 900 2408 902 2417
rect 1676 2382 1728 2388
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 846 2343 902 2352
rect 1688 1193 1716 2382
rect 8024 2304 8076 2310
rect 8392 2304 8444 2310
rect 8024 2246 8076 2252
rect 8390 2272 8392 2281
rect 8444 2272 8446 2281
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 8036 1193 8064 2246
rect 8390 2207 8446 2216
rect 1674 1184 1730 1193
rect 1674 1119 1730 1128
rect 8022 1184 8078 1193
rect 8022 1119 8078 1128
<< via2 >>
rect 1490 8744 1546 8800
rect 8022 8744 8078 8800
rect 846 7520 902 7576
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 8390 7656 8446 7712
rect 938 6568 994 6624
rect 1398 5480 1454 5536
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 846 4564 848 4584
rect 848 4564 900 4584
rect 900 4564 902 4584
rect 846 4528 902 4564
rect 846 3476 848 3496
rect 848 3476 900 3496
rect 900 3476 902 3496
rect 846 3440 902 3476
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 8390 6604 8392 6624
rect 8392 6604 8444 6624
rect 8444 6604 8446 6624
rect 8390 6568 8446 6604
rect 8206 5516 8208 5536
rect 8208 5516 8260 5536
rect 8260 5516 8262 5536
rect 8206 5480 8262 5516
rect 8390 4428 8392 4448
rect 8392 4428 8444 4448
rect 8444 4428 8446 4448
rect 8390 4392 8446 4428
rect 8390 3340 8392 3360
rect 8392 3340 8444 3360
rect 8444 3340 8446 3360
rect 8390 3304 8446 3340
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 8390 2252 8392 2272
rect 8392 2252 8444 2272
rect 8444 2252 8446 2272
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 8390 2216 8446 2252
rect 1674 1128 1730 1184
rect 8022 1128 8078 1184
<< metal3 >>
rect 0 8802 800 8832
rect 1485 8802 1551 8805
rect 0 8800 1551 8802
rect 0 8744 1490 8800
rect 1546 8744 1551 8800
rect 0 8742 1551 8744
rect 0 8712 800 8742
rect 1485 8739 1551 8742
rect 8017 8802 8083 8805
rect 9200 8802 10000 8832
rect 8017 8800 10000 8802
rect 8017 8744 8022 8800
rect 8078 8744 10000 8800
rect 8017 8742 10000 8744
rect 8017 8739 8083 8742
rect 9200 8712 10000 8742
rect 0 7714 800 7744
rect 8385 7714 8451 7717
rect 9200 7714 10000 7744
rect 0 7624 858 7714
rect 8385 7712 10000 7714
rect 8385 7656 8390 7712
rect 8446 7656 10000 7712
rect 8385 7654 10000 7656
rect 8385 7651 8451 7654
rect 798 7581 858 7624
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 9200 7624 10000 7654
rect 7606 7583 7922 7584
rect 798 7576 907 7581
rect 798 7520 846 7576
rect 902 7520 907 7576
rect 798 7518 907 7520
rect 841 7515 907 7518
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 0 6626 800 6656
rect 933 6626 999 6629
rect 0 6624 999 6626
rect 0 6568 938 6624
rect 994 6568 999 6624
rect 0 6566 999 6568
rect 0 6536 800 6566
rect 933 6563 999 6566
rect 8385 6626 8451 6629
rect 9200 6626 10000 6656
rect 8385 6624 10000 6626
rect 8385 6568 8390 6624
rect 8446 6568 10000 6624
rect 8385 6566 10000 6568
rect 8385 6563 8451 6566
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 9200 6536 10000 6566
rect 7606 6495 7922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 8201 5538 8267 5541
rect 9200 5538 10000 5568
rect 8201 5536 10000 5538
rect 8201 5480 8206 5536
rect 8262 5480 10000 5536
rect 8201 5478 10000 5480
rect 8201 5475 8267 5478
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 9200 5448 10000 5478
rect 7606 5407 7922 5408
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 841 4586 907 4589
rect 798 4584 907 4586
rect 798 4528 846 4584
rect 902 4528 907 4584
rect 798 4523 907 4528
rect 798 4480 858 4523
rect 0 4390 858 4480
rect 8385 4450 8451 4453
rect 9200 4450 10000 4480
rect 8385 4448 10000 4450
rect 8385 4392 8390 4448
rect 8446 4392 10000 4448
rect 8385 4390 10000 4392
rect 0 4360 800 4390
rect 8385 4387 8451 4390
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 9200 4360 10000 4390
rect 7606 4319 7922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 841 3498 907 3501
rect 798 3496 907 3498
rect 798 3440 846 3496
rect 902 3440 907 3496
rect 798 3435 907 3440
rect 798 3392 858 3435
rect 0 3302 858 3392
rect 8385 3362 8451 3365
rect 9200 3362 10000 3392
rect 8385 3360 10000 3362
rect 8385 3304 8390 3360
rect 8446 3304 10000 3360
rect 8385 3302 10000 3304
rect 0 3272 800 3302
rect 8385 3299 8451 3302
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 9200 3272 10000 3302
rect 7606 3231 7922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 841 2410 907 2413
rect 798 2408 907 2410
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2347 907 2352
rect 798 2304 858 2347
rect 0 2214 858 2304
rect 8385 2274 8451 2277
rect 9200 2274 10000 2304
rect 8385 2272 10000 2274
rect 8385 2216 8390 2272
rect 8446 2216 10000 2272
rect 8385 2214 10000 2216
rect 0 2184 800 2214
rect 8385 2211 8451 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 9200 2184 10000 2214
rect 7606 2143 7922 2144
rect 0 1186 800 1216
rect 1669 1186 1735 1189
rect 0 1184 1735 1186
rect 0 1128 1674 1184
rect 1730 1128 1735 1184
rect 0 1126 1735 1128
rect 0 1096 800 1126
rect 1669 1123 1735 1126
rect 8017 1186 8083 1189
rect 9200 1186 10000 1216
rect 8017 1184 10000 1186
rect 8017 1128 8022 1184
rect 8078 1128 10000 1184
rect 8017 1126 10000 1128
rect 8017 1123 8083 1126
rect 9200 1096 10000 1126
<< via3 >>
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
<< metal4 >>
rect 1944 7104 2264 7664
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 7648 2924 7664
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 7104 7264 7664
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 7648 7924 7664
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
<< via4 >>
rect 1986 3058 2222 3294
rect 2646 3718 2882 3954
rect 6986 3058 7222 3294
rect 7646 3718 7882 3954
<< metal5 >>
rect 1056 3954 8880 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 8880 3954
rect 1056 3676 8880 3718
rect 1056 3294 8880 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 8880 3294
rect 1056 3016 8880 3058
use sky130_fd_sc_hd__or4_2  _09_
timestamp 0
transform -1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _10_
timestamp 0
transform -1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _11_
timestamp 0
transform 1 0 1932 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _12_
timestamp 0
transform -1 0 7452 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _13_
timestamp 0
transform 1 0 5244 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _14_
timestamp 0
transform -1 0 2484 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _15_
timestamp 0
transform 1 0 2392 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _16_
timestamp 0
transform -1 0 6256 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 0
transform -1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _18_
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _19_
timestamp 0
transform 1 0 7268 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _20_
timestamp 0
transform 1 0 2208 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _21_
timestamp 0
transform -1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 0
transform 1 0 6072 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 0
transform -1 0 6716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _24_
timestamp 0
transform -1 0 6992 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 0
transform -1 0 5060 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_11
timestamp 0
transform 1 0 2116 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_17
timestamp 0
transform 1 0 2668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_29
timestamp 0
transform 1 0 3772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_37
timestamp 0
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_43
timestamp 0
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_6
timestamp 0
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_18
timestamp 0
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 0
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_49
timestamp 0
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_60
timestamp 0
transform 1 0 6624 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_72
timestamp 0
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_76
timestamp 0
transform 1 0 8096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_7
timestamp 0
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 0
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 0
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 0
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_36
timestamp 0
transform 1 0 4416 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_48
timestamp 0
transform 1 0 5520 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_60
timestamp 0
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_72
timestamp 0
transform 1 0 7728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_76
timestamp 0
transform 1 0 8096 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_11
timestamp 0
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_20
timestamp 0
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_32
timestamp 0
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_44
timestamp 0
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_61
timestamp 0
transform 1 0 6716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_73
timestamp 0
transform 1 0 7820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_6
timestamp 0
transform 1 0 1656 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_52
timestamp 0
transform 1 0 5888 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_64
timestamp 0
transform 1 0 6992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_74
timestamp 0
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_14
timestamp 0
transform 1 0 2392 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_26
timestamp 0
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_38
timestamp 0
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_50
timestamp 0
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_64
timestamp 0
transform 1 0 6992 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_76
timestamp 0
transform 1 0 8096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_80
timestamp 0
transform 1 0 8464 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_13
timestamp 0
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 0
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_59
timestamp 0
transform 1 0 6532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_69
timestamp 0
transform 1 0 7452 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_13
timestamp 0
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_25
timestamp 0
transform 1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_36
timestamp 0
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_48
timestamp 0
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform 1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_22
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_23
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_24
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_25
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_26
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_27
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_28
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_29
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_30
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_31
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
<< labels >>
rlabel metal1 s 4968 7616 4968 7616 4 VGND
rlabel metal1 s 4968 7072 4968 7072 4 VPWR
rlabel metal2 s 3910 5508 3910 5508 4 _00_
rlabel metal1 s 5382 5780 5382 5780 4 _01_
rlabel metal2 s 7406 6596 7406 6596 4 _02_
rlabel metal2 s 6210 3740 6210 3740 4 _03_
rlabel metal1 s 3266 4998 3266 4998 4 _04_
rlabel metal2 s 5750 5236 5750 5236 4 _05_
rlabel metal1 s 6302 6290 6302 6290 4 _06_
rlabel metal1 s 6348 3706 6348 3706 4 _07_
rlabel metal2 s 6486 5916 6486 5916 4 _08_
rlabel metal3 s 1096 8772 1096 8772 4 in[0]
rlabel metal3 s 0 7624 800 7744 4 in[1]
port 4 nsew
rlabel metal3 s 820 6596 820 6596 4 in[2]
rlabel metal3 s 1050 5508 1050 5508 4 in[3]
rlabel metal3 s 0 4360 800 4480 4 in[4]
port 7 nsew
rlabel metal3 s 0 3272 800 3392 4 in[5]
port 8 nsew
rlabel metal3 s 0 2184 800 2304 4 in[6]
port 9 nsew
rlabel metal3 s 1188 1156 1188 1156 4 in[7]
rlabel metal1 s 1978 3026 1978 3026 4 net1
rlabel metal1 s 8050 5882 8050 5882 4 net10
rlabel metal2 s 7498 6052 7498 6052 4 net11
rlabel metal2 s 7590 5882 7590 5882 4 net12
rlabel metal1 s 7774 4590 7774 4590 4 net13
rlabel metal2 s 6670 4522 6670 4522 4 net14
rlabel metal1 s 2254 6664 2254 6664 4 net15
rlabel metal2 s 4370 4794 4370 4794 4 net16
rlabel metal1 s 1886 2822 1886 2822 4 net2
rlabel metal2 s 4186 4386 4186 4386 4 net3
rlabel metal2 s 4094 5474 4094 5474 4 net4
rlabel metal1 s 2300 5678 2300 5678 4 net5
rlabel metal2 s 2530 5338 2530 5338 4 net6
rlabel metal1 s 1794 4114 1794 4114 4 net7
rlabel metal1 s 2944 2618 2944 2618 4 net8
rlabel metal1 s 6532 2890 6532 2890 4 net9
rlabel metal2 s 8050 8143 8050 8143 4 out[0]
rlabel metal2 s 8418 7599 8418 7599 4 out[1]
rlabel metal3 s 8418 6613 8418 6613 4 out[2]
rlabel metal1 s 8326 5542 8326 5542 4 out[3]
rlabel metal3 s 8418 4437 8418 4437 4 out[4]
rlabel metal3 s 8418 3349 8418 3349 4 out[5]
rlabel metal3 s 8418 2261 8418 2261 4 out[6]
rlabel metal2 s 8050 1717 8050 1717 4 out[7]
flabel metal5 s 1056 3676 8880 3996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 7604 2128 7924 7664 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2604 2128 2924 7664 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3016 8880 3336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 6944 2128 7264 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1944 2128 2264 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 8712 800 8832 0 FreeSans 600 0 0 0 in[0]
port 3 nsew
flabel metal3 s 400 7684 400 7684 0 FreeSans 600 0 0 0 in[1]
flabel metal3 s 0 6536 800 6656 0 FreeSans 600 0 0 0 in[2]
port 5 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 in[3]
port 6 nsew
flabel metal3 s 400 4420 400 4420 0 FreeSans 600 0 0 0 in[4]
flabel metal3 s 400 3332 400 3332 0 FreeSans 600 0 0 0 in[5]
flabel metal3 s 400 2244 400 2244 0 FreeSans 600 0 0 0 in[6]
flabel metal3 s 0 1096 800 1216 0 FreeSans 600 0 0 0 in[7]
port 10 nsew
flabel metal3 s 9200 8712 10000 8832 0 FreeSans 600 0 0 0 out[0]
port 11 nsew
flabel metal3 s 9200 7624 10000 7744 0 FreeSans 600 0 0 0 out[1]
port 12 nsew
flabel metal3 s 9200 6536 10000 6656 0 FreeSans 600 0 0 0 out[2]
port 13 nsew
flabel metal3 s 9200 5448 10000 5568 0 FreeSans 600 0 0 0 out[3]
port 14 nsew
flabel metal3 s 9200 4360 10000 4480 0 FreeSans 600 0 0 0 out[4]
port 15 nsew
flabel metal3 s 9200 3272 10000 3392 0 FreeSans 600 0 0 0 out[5]
port 16 nsew
flabel metal3 s 9200 2184 10000 2304 0 FreeSans 600 0 0 0 out[6]
port 17 nsew
flabel metal3 s 9200 1096 10000 1216 0 FreeSans 600 0 0 0 out[7]
port 18 nsew
<< properties >>
string FIXED_BBOX 0 0 10000 10000
<< end >>
